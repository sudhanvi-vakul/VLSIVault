class alu_smoke_test extends uvm_test;
  `uvm_component_utils(alu_smoke_test);
  
  alu_env env;
  
  function new(string name = "alu_smoke_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = alu_env::type_id::create("env", this);
  endfunction
  
  virtual task run_phase(uvm_phase phase);
    
    alu_directed_seq seq;
    
    phase.raise_objection(this);

    seq = alu_directed_seq::type_id::create("seq");
    seq.start(env.agent.seqr);
    #500;
    phase.drop_objection(this);
    
  endtask
endclass
    