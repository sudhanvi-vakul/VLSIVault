class alu_env extends uvm_env;
  `uvm_component_utils(alu_env)
  
  alu_agent agent;
  alu_scoreboard scoreboard;
  
  function new(string name = "alu_env", uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("ENV", "In build_phase", UVM_LOW)
    agent = alu_agent::type_id::create("agent", this);
    scoreboard = alu_scoreboard::type_id::create("scoreboard", this);
  endfunction
  
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    `uvm_info("ENV", "In connect_phase", UVM_LOW)
    agent.mon.ap.connect(scoreboard.imp);
  endfunction
  
endclass