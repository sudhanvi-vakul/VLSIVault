`include "uvm_macros.svh"
module uvm_smoke;
  import uvm_pkg::*;
  initial begin
    `uvm_info("UVM_SMOKE", "UVM is available", UVM_LOW)
  end
endmodule

